library ieee;
use ieee.std_logic_1164.all;

entity enpulsare is
	port(clk, reset : in std_logic; -- reset is active high.
	     x : in std_logic; -- x
	     u : out std_logic);
end entity;

architecture behav of enpulsare is
begin
end architecture;

