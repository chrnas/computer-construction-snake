library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity CHAR_ROM is
    port(
      CR_addr       : in unsigned (9 downto 0);
      vgaRed        : out std_logic_vector(2 downto 0);
      vgaGreen      : out std_logic_vector(2 downto 0);
      vgaBlue       : out std_logic_vector(2 downto 1));
  end CHAR_ROM;

architecture Behavioral of CHAR_ROM is

type ch_mem_t is array (0 to 600) of unsigned(2 downto 0);
constant ch_mem_c : ch_mem_t :=
  (
    -- Border   (x"0")
    "111", "111", "111", "111", "111", "111", "111", "111",
    "111", "111", "111", "111", "111", "111", "111", "111",
    "111", "111", "111", "111", "111", "111", "111", "111",
    "111", "111", "111", "111", "111", "111", "111", "111",
    "111", "111", "111", "111", "111", "111", "111", "111",
    "111", "111", "111", "111", "111", "111", "111", "111",
    "111", "111", "111", "111", "111", "111", "111", "111",
    "111", "111", "111", "111", "111", "111", "111", "111",

    -- Background   (x"1")
    "111", "000", "000", "000", "000", "000", "000", "111",
    "000", "000", "000", "000", "000", "000", "000", "000",
    "000", "000", "000", "000", "000", "000", "000", "000",
    "000", "000", "000", "000", "000", "000", "000", "000",
    "000", "000", "000", "000", "000", "000", "000", "000",
    "000", "000", "000", "000", "000", "000", "000", "000",
    "000", "000", "000", "000", "000", "000", "000", "000",
    "111", "000", "000", "000", "000", "000", "000", "111",

    -- Apple   (x"2")
    "000", "000", "100", "100", "100", "100", "000", "000",
    "000", "100", "100", "100", "100", "100", "100", "000",
    "100", "100", "100", "100", "100", "100", "100", "100",
    "100", "100", "100", "100", "100", "100", "100", "100",
    "100", "100", "100", "100", "100", "100", "100", "100",
    "100", "100", "100", "100", "100", "100", "100", "100",
    "000", "100", "100", "100", "100", "100", "100", "000",
    "000", "000", "100", "100", "100", "100", "000", "000",

    -- Snake Up   (x"3")
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "000",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",

    -- Snake Down   (x"4")
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "000",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",

    -- Snake Left    (x"5")
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "000",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",

    -- Snake Right   (x"6")
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "000",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",
    "010", "010", "010", "010", "010", "010", "010", "010",

    others => (others => '0')
  );

  signal ch_mem : ch_mem_t := ch_mem_c;

  signal temp : unsigned(9 downto 0);

  begin

    temp <= CR_addr;

    --type code for outputs
    vgaRed(0) <= ch_mem(to_integer(temp))(2);
    vgaRed(1) <= ch_mem(to_integer(temp))(2);
    vgaRed(2) <= ch_mem(to_integer(temp))(2);
    vgaGreen(0) <= ch_mem(to_integer(temp))(1);
    vgaGreen(1) <= ch_mem(to_integer(temp))(1);
    vgaGreen(2) <= ch_mem(to_integer(temp))(1);
    vgaBlue(1) <= ch_mem(to_integer(temp))(0);
    vgaBlue(2) <= ch_mem(to_integer(temp))(0);

  end Behavioral;
